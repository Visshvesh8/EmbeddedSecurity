module _xor(a, b, op);
    input a,b;
    output op;
    
    assign op = a^b;

endmodule